# SCHISM sflux input file (sflux_rad_*.nc)
# Based on NARR file format: http://ccrm.vims.edu/yinglong/wiki_files/NARR/

netcdf sflux_rad {
dimensions:
	nx_grid = 0 ;
	ny_grid = 0 ;
	time = 0 ; 
variables:
	float time(time) ;
		time:long_name = "Time" ;
		time:standard_name = "time" ;
		time:units = "seconds since XXXX" ;
		time:base_date = XXXX ;
	float lon(ny_grid, nx_grid) ;
		lon:long_name = "Longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	float lat(ny_grid, nx_grid) ;
		lat:long_name = "Latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	float dlwrf(time, ny_grid, nx_grid) ;
		dlwrf:long_name = "Downward Long Wave Radiation Flux" ;
		dlwrf:standard_name = "surface_downwelling_longwave_flux_in_air" ;
		dlwrf:units = "W/m^2" ;
	float dswrf(time, ny_grid, nx_grid) ;
		dswrf:long_name = "Downward Short Wave Radiation Flux" ;
		dswrf:standard_name = "surface_downwelling_shortwave_flux_in_air" ;
		dswrf:units = "W/m^2" ;

// global attributes:
        :type = "" ;
        :title = "" ;
        :Conventions = "CF-1.0" ;
}