# SCHISM hotstart file (hotstart.nc)

netcdf hotstart {
dimensions:
        node = 77051 ;
        elem = 145682 ;
        side = 222751 ;
        nVert = 11 ;
        ntracers = 2 ;
        one = 1 ;
        three = 3 ;
        two = 2 ;
        four = 4 ;
        five = 5 ;
        six = 6 ;
        seven = 7 ;
        eight = 8 ;
        nine = 9 ;
        one_new = 1 ;
variables:
        double time(one_new) ;
                time:long_name = "" ;
                time:units = "" ;
                time:time = "" ;
                time:_FillValue = 1.e+20 ;
        int iths(one_new) ;
                iths:long_name = "iteration number" ;
                iths:units = "" ;
                iths:time = "" ;
                iths:_FillValue = 1.e+20 ;
        int ifile(one_new) ;
                ifile:long_name = "file number" ;
                ifile:units = "" ;
                ifile:time = "" ;
                ifile:_FillValue = 1.e+20 ;
        int idry_e(elem) ;
                idry_e:long_name = "wet/dry flag at elements" ;
                idry_e:units = "" ;
                idry_e:time = "" ;
                idry_e:_FillValue = 1.e+20 ;
        int idry_s(side) ;
                idry_s:long_name = "wet/dry flag at sides" ;
                idry_s:units = "" ;
                idry_s:time = "" ;
                idry_s:_FillValue = 1.e+20 ;
        int idry(node) ;
                idry:long_name = "wet/dry flag at nodes" ;
                idry:units = "" ;
                idry:time = "" ;
                idry:_FillValue = 1.e+20 ;
        double eta2(node) ;
                eta2:long_name = "elevation at nodes at current timestep" ;
                eta2:units = "" ;
                eta2:time = "" ;
                eta2:_FillValue = 1.e+20 ;
        double su2(side, nVert) ;
                su2:long_name = "u-velocity at side centers" ;
                su2:units = "" ;
                su2:time = "" ;
                su2:_FillValue = 1.e+20 ;
        double sv2(side, nVert) ;
                sv2:long_name = "v-velocity at side centers" ;
                sv2:units = "" ;
                sv2:time = "" ;
                sv2:_FillValue = 1.e+20 ;
        double we(elem, nVert) ;
                we:long_name = "vertical velocity at element centers, calculated using F.V.M." ;
                we:units = "" ;
                we:time = "" ;
                we:_FillValue = 1.e+20 ;
        double tr_el(elem, nVert, ntracers) ;
                tr_el:long_name = "tracer concentration at elements" ;
                tr_el:units = "" ;
                tr_el:time = "" ;
                tr_el:_FillValue = 1.e+20 ;
        double tr_nd0(node, nVert, ntracers) ;
                tr_nd0:long_name = "initial tracer concentration at nodes" ;
                tr_nd0:units = "" ;
                tr_nd0:time = "" ;
                tr_nd0:_FillValue = 1.e+20 ;
        double tr_nd(node, nVert, ntracers) ;
                tr_nd:long_name = "tracer concentration at nodes" ;
                tr_nd:units = "" ;
                tr_nd:time = "" ;
                tr_nd:_FillValue = 1.e+20 ;
        double q2(node, nVert) ;
                q2:long_name = "turbulent kinetic energy at sides and half levels" ;
                q2:units = "" ;
                q2:time = "" ;
                q2:_FillValue = 1.e+20 ;
        double xl(node, nVert) ;
                xl:long_name = "turbulent mixing length at sides and half levels" ;
                xl:units = "" ;
                xl:time = "" ;
                xl:_FillValue = 1.e+20 ;
        double dfv(node, nVert) ;
                dfv:long_name = "viscosity at nodes" ;
                dfv:units = "" ;
                dfv:time = "" ;
                dfv:_FillValue = 1.e+20 ;
        double dfh(node, nVert) ;
                dfh:long_name = "diffusivity at nodes" ;
                dfh:units = "" ;
                dfh:time = "" ;
                dfh:_FillValue = 1.e+20 ;
        double dfq1(node, nVert) ;
                dfq1:long_name = "diffmin" ;
                dfq1:units = "" ;
                dfq1:time = "" ;
                dfq1:_FillValue = 1.e+20 ;
        double dfq2(node, nVert) ;
                dfq2:long_name = "diffmax" ;
                dfq2:units = "" ;
                dfq2:time = "" ;
                dfq2:_FillValue = 1.e+20 ;
// global attributes:
        :type = "" ;
        :title = "" ;
}